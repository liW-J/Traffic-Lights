-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Mon Nov 30 20:47:42 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY traffic IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		EN :  IN  STD_LOGIC;
		RST :  IN  STD_LOGIC;
		DX1 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		DX2 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		LIGHT :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		LIGHTA :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		NB1 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		NB2 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END traffic;

ARCHITECTURE bdf_type OF traffic IS 

COMPONENT control
	PORT(CLK : IN STD_LOGIC;
		 EN : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 DX : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 NB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT display
	PORT(S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 LIGHT : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 LIGHTA : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT time
	PORT(CLK : IN STD_LOGIC;
		 RST : IN STD_LOGIC;
		 EN : IN STD_LOGIC;
		 S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 DX7 : OUT STD_LOGIC;
		 DX6 : OUT STD_LOGIC;
		 DX5 : OUT STD_LOGIC;
		 DX4 : OUT STD_LOGIC;
		 DX3 : OUT STD_LOGIC;
		 DX2 : OUT STD_LOGIC;
		 DX1 : OUT STD_LOGIC;
		 DX0 : OUT STD_LOGIC;
		 DX13 : OUT STD_LOGIC;
		 DX12 : OUT STD_LOGIC;
		 DX11 : OUT STD_LOGIC;
		 DX10 : OUT STD_LOGIC;
		 DX23 : OUT STD_LOGIC;
		 DX22 : OUT STD_LOGIC;
		 DX21 : OUT STD_LOGIC;
		 DX20 : OUT STD_LOGIC;
		 NB7 : OUT STD_LOGIC;
		 NB6 : OUT STD_LOGIC;
		 NB5 : OUT STD_LOGIC;
		 NB4 : OUT STD_LOGIC;
		 NB3 : OUT STD_LOGIC;
		 NB2 : OUT STD_LOGIC;
		 NB1 : OUT STD_LOGIC;
		 NB0 : OUT STD_LOGIC;
		 NB13 : OUT STD_LOGIC;
		 NB12 : OUT STD_LOGIC;
		 NB11 : OUT STD_LOGIC;
		 NB10 : OUT STD_LOGIC;
		 NB23 : OUT STD_LOGIC;
		 NB22 : OUT STD_LOGIC;
		 NB21 : OUT STD_LOGIC;
		 NB20 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL	GDFX_TEMP_SIGNAL_30 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_31 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_32 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_33 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_26 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_27 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_28 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_29 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_18 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_19 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_20 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_21 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_22 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_23 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_24 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_25 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_14 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_15 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_16 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_17 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_10 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_11 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_12 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_13 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_8 :  STD_LOGIC;
SIGNAL	GDFX_TEMP_SIGNAL_9 :  STD_LOGIC;

BEGIN 

NB23 <= GDFX_TEMP_SIGNAL_30;
NB22 <= GDFX_TEMP_SIGNAL_30;
NB21 <= GDFX_TEMP_SIGNAL_30;
NB20 <= GDFX_TEMP_SIGNAL_30;

NB23 <= GDFX_TEMP_SIGNAL_31;
NB22 <= GDFX_TEMP_SIGNAL_31;
NB21 <= GDFX_TEMP_SIGNAL_31;
NB20 <= GDFX_TEMP_SIGNAL_31;

NB23 <= GDFX_TEMP_SIGNAL_32;
NB22 <= GDFX_TEMP_SIGNAL_32;
NB21 <= GDFX_TEMP_SIGNAL_32;
NB20 <= GDFX_TEMP_SIGNAL_32;

NB23 <= GDFX_TEMP_SIGNAL_33;
NB22 <= GDFX_TEMP_SIGNAL_33;
NB21 <= GDFX_TEMP_SIGNAL_33;
NB20 <= GDFX_TEMP_SIGNAL_33;

NB13 <= GDFX_TEMP_SIGNAL_26;
NB12 <= GDFX_TEMP_SIGNAL_26;
NB11 <= GDFX_TEMP_SIGNAL_26;
NB10 <= GDFX_TEMP_SIGNAL_26;

NB13 <= GDFX_TEMP_SIGNAL_27;
NB12 <= GDFX_TEMP_SIGNAL_27;
NB11 <= GDFX_TEMP_SIGNAL_27;
NB10 <= GDFX_TEMP_SIGNAL_27;

NB13 <= GDFX_TEMP_SIGNAL_28;
NB12 <= GDFX_TEMP_SIGNAL_28;
NB11 <= GDFX_TEMP_SIGNAL_28;
NB10 <= GDFX_TEMP_SIGNAL_28;

NB13 <= GDFX_TEMP_SIGNAL_29;
NB12 <= GDFX_TEMP_SIGNAL_29;
NB11 <= GDFX_TEMP_SIGNAL_29;
NB10 <= GDFX_TEMP_SIGNAL_29;

GDFX_TEMP_SIGNAL_1 <= (NB7 & NB6 & NB5 & NB4 & NB3 & NB2 & NB1 & NB0);
NB7 <= GDFX_TEMP_SIGNAL_18;
NB6 <= GDFX_TEMP_SIGNAL_18;
NB5 <= GDFX_TEMP_SIGNAL_18;
NB4 <= GDFX_TEMP_SIGNAL_18;
NB3 <= GDFX_TEMP_SIGNAL_18;
NB2 <= GDFX_TEMP_SIGNAL_18;
NB1 <= GDFX_TEMP_SIGNAL_18;
NB0 <= GDFX_TEMP_SIGNAL_18;

NB7 <= GDFX_TEMP_SIGNAL_19;
NB6 <= GDFX_TEMP_SIGNAL_19;
NB5 <= GDFX_TEMP_SIGNAL_19;
NB4 <= GDFX_TEMP_SIGNAL_19;
NB3 <= GDFX_TEMP_SIGNAL_19;
NB2 <= GDFX_TEMP_SIGNAL_19;
NB1 <= GDFX_TEMP_SIGNAL_19;
NB0 <= GDFX_TEMP_SIGNAL_19;

NB7 <= GDFX_TEMP_SIGNAL_20;
NB6 <= GDFX_TEMP_SIGNAL_20;
NB5 <= GDFX_TEMP_SIGNAL_20;
NB4 <= GDFX_TEMP_SIGNAL_20;
NB3 <= GDFX_TEMP_SIGNAL_20;
NB2 <= GDFX_TEMP_SIGNAL_20;
NB1 <= GDFX_TEMP_SIGNAL_20;
NB0 <= GDFX_TEMP_SIGNAL_20;

NB7 <= GDFX_TEMP_SIGNAL_21;
NB6 <= GDFX_TEMP_SIGNAL_21;
NB5 <= GDFX_TEMP_SIGNAL_21;
NB4 <= GDFX_TEMP_SIGNAL_21;
NB3 <= GDFX_TEMP_SIGNAL_21;
NB2 <= GDFX_TEMP_SIGNAL_21;
NB1 <= GDFX_TEMP_SIGNAL_21;
NB0 <= GDFX_TEMP_SIGNAL_21;

NB7 <= GDFX_TEMP_SIGNAL_22;
NB6 <= GDFX_TEMP_SIGNAL_22;
NB5 <= GDFX_TEMP_SIGNAL_22;
NB4 <= GDFX_TEMP_SIGNAL_22;
NB3 <= GDFX_TEMP_SIGNAL_22;
NB2 <= GDFX_TEMP_SIGNAL_22;
NB1 <= GDFX_TEMP_SIGNAL_22;
NB0 <= GDFX_TEMP_SIGNAL_22;

NB7 <= GDFX_TEMP_SIGNAL_23;
NB6 <= GDFX_TEMP_SIGNAL_23;
NB5 <= GDFX_TEMP_SIGNAL_23;
NB4 <= GDFX_TEMP_SIGNAL_23;
NB3 <= GDFX_TEMP_SIGNAL_23;
NB2 <= GDFX_TEMP_SIGNAL_23;
NB1 <= GDFX_TEMP_SIGNAL_23;
NB0 <= GDFX_TEMP_SIGNAL_23;

NB7 <= GDFX_TEMP_SIGNAL_24;
NB6 <= GDFX_TEMP_SIGNAL_24;
NB5 <= GDFX_TEMP_SIGNAL_24;
NB4 <= GDFX_TEMP_SIGNAL_24;
NB3 <= GDFX_TEMP_SIGNAL_24;
NB2 <= GDFX_TEMP_SIGNAL_24;
NB1 <= GDFX_TEMP_SIGNAL_24;
NB0 <= GDFX_TEMP_SIGNAL_24;

NB7 <= GDFX_TEMP_SIGNAL_25;
NB6 <= GDFX_TEMP_SIGNAL_25;
NB5 <= GDFX_TEMP_SIGNAL_25;
NB4 <= GDFX_TEMP_SIGNAL_25;
NB3 <= GDFX_TEMP_SIGNAL_25;
NB2 <= GDFX_TEMP_SIGNAL_25;
NB1 <= GDFX_TEMP_SIGNAL_25;
NB0 <= GDFX_TEMP_SIGNAL_25;

DX23 <= GDFX_TEMP_SIGNAL_14;
DX22 <= GDFX_TEMP_SIGNAL_14;
DX21 <= GDFX_TEMP_SIGNAL_14;
DX20 <= GDFX_TEMP_SIGNAL_14;

DX23 <= GDFX_TEMP_SIGNAL_15;
DX22 <= GDFX_TEMP_SIGNAL_15;
DX21 <= GDFX_TEMP_SIGNAL_15;
DX20 <= GDFX_TEMP_SIGNAL_15;

DX23 <= GDFX_TEMP_SIGNAL_16;
DX22 <= GDFX_TEMP_SIGNAL_16;
DX21 <= GDFX_TEMP_SIGNAL_16;
DX20 <= GDFX_TEMP_SIGNAL_16;

DX23 <= GDFX_TEMP_SIGNAL_17;
DX22 <= GDFX_TEMP_SIGNAL_17;
DX21 <= GDFX_TEMP_SIGNAL_17;
DX20 <= GDFX_TEMP_SIGNAL_17;

DX13 <= GDFX_TEMP_SIGNAL_10;
DX12 <= GDFX_TEMP_SIGNAL_10;
DX11 <= GDFX_TEMP_SIGNAL_10;
DX10 <= GDFX_TEMP_SIGNAL_10;

DX13 <= GDFX_TEMP_SIGNAL_11;
DX12 <= GDFX_TEMP_SIGNAL_11;
DX11 <= GDFX_TEMP_SIGNAL_11;
DX10 <= GDFX_TEMP_SIGNAL_11;

DX13 <= GDFX_TEMP_SIGNAL_12;
DX12 <= GDFX_TEMP_SIGNAL_12;
DX11 <= GDFX_TEMP_SIGNAL_12;
DX10 <= GDFX_TEMP_SIGNAL_12;

DX13 <= GDFX_TEMP_SIGNAL_13;
DX12 <= GDFX_TEMP_SIGNAL_13;
DX11 <= GDFX_TEMP_SIGNAL_13;
DX10 <= GDFX_TEMP_SIGNAL_13;

GDFX_TEMP_SIGNAL_0 <= (DX7 & DX6 & DX5 & DX4 & DX3 & DX2 & DX1 & DX0);
DX7 <= GDFX_TEMP_SIGNAL_2;
DX6 <= GDFX_TEMP_SIGNAL_2;
DX5 <= GDFX_TEMP_SIGNAL_2;
DX4 <= GDFX_TEMP_SIGNAL_2;
DX3 <= GDFX_TEMP_SIGNAL_2;
DX2 <= GDFX_TEMP_SIGNAL_2;
DX1 <= GDFX_TEMP_SIGNAL_2;
DX0 <= GDFX_TEMP_SIGNAL_2;

DX7 <= GDFX_TEMP_SIGNAL_3;
DX6 <= GDFX_TEMP_SIGNAL_3;
DX5 <= GDFX_TEMP_SIGNAL_3;
DX4 <= GDFX_TEMP_SIGNAL_3;
DX3 <= GDFX_TEMP_SIGNAL_3;
DX2 <= GDFX_TEMP_SIGNAL_3;
DX1 <= GDFX_TEMP_SIGNAL_3;
DX0 <= GDFX_TEMP_SIGNAL_3;

DX7 <= GDFX_TEMP_SIGNAL_4;
DX6 <= GDFX_TEMP_SIGNAL_4;
DX5 <= GDFX_TEMP_SIGNAL_4;
DX4 <= GDFX_TEMP_SIGNAL_4;
DX3 <= GDFX_TEMP_SIGNAL_4;
DX2 <= GDFX_TEMP_SIGNAL_4;
DX1 <= GDFX_TEMP_SIGNAL_4;
DX0 <= GDFX_TEMP_SIGNAL_4;

DX7 <= GDFX_TEMP_SIGNAL_5;
DX6 <= GDFX_TEMP_SIGNAL_5;
DX5 <= GDFX_TEMP_SIGNAL_5;
DX4 <= GDFX_TEMP_SIGNAL_5;
DX3 <= GDFX_TEMP_SIGNAL_5;
DX2 <= GDFX_TEMP_SIGNAL_5;
DX1 <= GDFX_TEMP_SIGNAL_5;
DX0 <= GDFX_TEMP_SIGNAL_5;

DX7 <= GDFX_TEMP_SIGNAL_6;
DX6 <= GDFX_TEMP_SIGNAL_6;
DX5 <= GDFX_TEMP_SIGNAL_6;
DX4 <= GDFX_TEMP_SIGNAL_6;
DX3 <= GDFX_TEMP_SIGNAL_6;
DX2 <= GDFX_TEMP_SIGNAL_6;
DX1 <= GDFX_TEMP_SIGNAL_6;
DX0 <= GDFX_TEMP_SIGNAL_6;

DX7 <= GDFX_TEMP_SIGNAL_7;
DX6 <= GDFX_TEMP_SIGNAL_7;
DX5 <= GDFX_TEMP_SIGNAL_7;
DX4 <= GDFX_TEMP_SIGNAL_7;
DX3 <= GDFX_TEMP_SIGNAL_7;
DX2 <= GDFX_TEMP_SIGNAL_7;
DX1 <= GDFX_TEMP_SIGNAL_7;
DX0 <= GDFX_TEMP_SIGNAL_7;

DX7 <= GDFX_TEMP_SIGNAL_8;
DX6 <= GDFX_TEMP_SIGNAL_8;
DX5 <= GDFX_TEMP_SIGNAL_8;
DX4 <= GDFX_TEMP_SIGNAL_8;
DX3 <= GDFX_TEMP_SIGNAL_8;
DX2 <= GDFX_TEMP_SIGNAL_8;
DX1 <= GDFX_TEMP_SIGNAL_8;
DX0 <= GDFX_TEMP_SIGNAL_8;

DX7 <= GDFX_TEMP_SIGNAL_9;
DX6 <= GDFX_TEMP_SIGNAL_9;
DX5 <= GDFX_TEMP_SIGNAL_9;
DX4 <= GDFX_TEMP_SIGNAL_9;
DX3 <= GDFX_TEMP_SIGNAL_9;
DX2 <= GDFX_TEMP_SIGNAL_9;
DX1 <= GDFX_TEMP_SIGNAL_9;
DX0 <= GDFX_TEMP_SIGNAL_9;



b2v_inst : control
PORT MAP(CLK => CLK,
		 EN => EN,
		 RST => RST,
		 DX => GDFX_TEMP_SIGNAL_0,
		 NB => GDFX_TEMP_SIGNAL_1,
		 Q => SYNTHESIZED_WIRE_2);


b2v_inst1 : display
PORT MAP(S => SYNTHESIZED_WIRE_2,
		 LIGHT => LIGHT,
		 LIGHTA => LIGHTA);


b2v_inst2 : time
PORT MAP(CLK => CLK,
		 RST => RST,
		 EN => EN,
		 S => SYNTHESIZED_WIRE_2,
		 DX7 => GDFX_TEMP_SIGNAL_2,
		 DX6 => GDFX_TEMP_SIGNAL_3,
		 DX5 => GDFX_TEMP_SIGNAL_4,
		 DX4 => GDFX_TEMP_SIGNAL_5,
		 DX3 => GDFX_TEMP_SIGNAL_6,
		 DX2 => GDFX_TEMP_SIGNAL_7,
		 DX1 => GDFX_TEMP_SIGNAL_8,
		 DX0 => GDFX_TEMP_SIGNAL_9,
		 DX13 => GDFX_TEMP_SIGNAL_10,
		 DX12 => GDFX_TEMP_SIGNAL_11,
		 DX11 => GDFX_TEMP_SIGNAL_12,
		 DX10 => GDFX_TEMP_SIGNAL_13,
		 DX23 => GDFX_TEMP_SIGNAL_14,
		 DX22 => GDFX_TEMP_SIGNAL_15,
		 DX21 => GDFX_TEMP_SIGNAL_16,
		 DX20 => GDFX_TEMP_SIGNAL_17,
		 NB7 => GDFX_TEMP_SIGNAL_18,
		 NB6 => GDFX_TEMP_SIGNAL_19,
		 NB5 => GDFX_TEMP_SIGNAL_20,
		 NB4 => GDFX_TEMP_SIGNAL_21,
		 NB3 => GDFX_TEMP_SIGNAL_22,
		 NB2 => GDFX_TEMP_SIGNAL_23,
		 NB1 => GDFX_TEMP_SIGNAL_24,
		 NB0 => GDFX_TEMP_SIGNAL_25,
		 NB13 => GDFX_TEMP_SIGNAL_26,
		 NB12 => GDFX_TEMP_SIGNAL_27,
		 NB11 => GDFX_TEMP_SIGNAL_28,
		 NB10 => GDFX_TEMP_SIGNAL_29,
		 NB23 => GDFX_TEMP_SIGNAL_30,
		 NB22 => GDFX_TEMP_SIGNAL_31,
		 NB21 => GDFX_TEMP_SIGNAL_32,
		 NB20 => GDFX_TEMP_SIGNAL_33);

DX1(3) <= DX13;
DX1(2) <= DX12;
DX1(1) <= DX11;
DX1(0) <= DX10;
DX2(3) <= DX23;
DX2(2) <= DX22;
DX2(1) <= DX21;
DX2(0) <= DX20;
NB1(3) <= NB13;
NB1(2) <= NB12;
NB1(1) <= NB11;
NB1(0) <= NB10;
NB2(3) <= NB23;
NB2(2) <= NB22;
NB2(1) <= NB21;
NB2(0) <= NB20;

END bdf_type;