library verilog;
use verilog.vl_types.all;
entity traffic_vlg_vec_tst is
end traffic_vlg_vec_tst;
