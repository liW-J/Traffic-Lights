LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY control IS
PORT(  CLK:IN STD_LOGIC;
       EN:IN STD_LOGIC;
       RST:IN STD_LOGIC;
       DX:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 NB:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 GLOBAL:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	    Q:OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		);
 END control;
 ARCHITECTURE behav OF control IS
 SIGNAL S:STD_LOGIC_VECTOR(1 DOWNTO 0):="11";
 SIGNAL COUNT: INTEGER RANGE 0 TO 15;
	 BEGIN

PROCESS (CLK,RST,EN)
BEGIN
    IF RST='0' THEN COUNT<=15;
	 ELSE IF RST='1' AND EN='0'THEN COUNT<=COUNT;
    ELSE
	 IF CLK'EVENT AND CLK='1' THEN
	 IF COUNT = 0 THEN COUNT<=15;
	 ELSE COUNT<=COUNT-1;
	 END IF;
	 END IF;
	 END IF;
	 END IF;
	 END PROCESS;
	 
PROCESS(CLK,COUNT,DX,NB,GLOBAL)
BEGIN
	IF GLOBAL="11" THEN
	IF CLK'EVENT AND CLK='0' AND COUNT= 15 THEN
			  IF(DX="00000001")OR(NB="00000001")THEN 
				S<=S+1; 				 			
			   ELSE S<=S;		   
			  END IF;
			 END IF;
	END IF;
	IF GLOBAL="01" THEN
		S<="00";
	END IF;
	IF GLOBAL="10" OR GLOBAL="00" THEN
		S<="10";
	END IF;
	Q<=S;
	END PROCESS;
	END behav;