-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "11/30/2020 16:14:46"
                                                            
-- Vhdl Test Bench template for design  :  control
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;                                               
USE ieee.std_logic_1164.all;                                

ENTITY control_vhd_tst IS
END control_vhd_tst;
ARCHITECTURE control_arch OF control_vhd_tst IS
-- constants
CONSTANT CLK_P : TIME := 31.25 ms;                                                 
-- signals                                                   
SIGNAL CLK : STD_LOGIC;
SIGNAL DX : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL EN : STD_LOGIC;
SIGNAL NB : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL Q : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL RST : STD_LOGIC;
COMPONENT control
	PORT (
	CLK : IN STD_LOGIC;
	DX : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	EN : IN STD_LOGIC;
	NB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	RST : IN STD_LOGIC
	);
END COMPONENT;
BEGIN
	i1 : control
	PORT MAP (
-- list connections between master ports and signals
	CLK => CLK,
	DX => DX,
	EN => EN,
	NB => NB,
	Q => Q,
	RST => RST
	);
init : PROCESS                                               
-- variable declarations                                     
BEGIN                                                        
        -- code that executes only once                      
WAIT;                                                       
END PROCESS init;                                           
always : PROCESS                                              
-- optional sensitivity list                                  
-- (        )                                                 
-- variable declarations                                      
BEGIN                                                         
  CLK <= '0';                   
  WAIT FOR CLK_P;
  CLK <= '1';
  WAIT FOR CLK_P;                                                         
END PROCESS always; 
RST <= '0', '1' AFTER 1*CLK_P;
EN <= '0', '1' AFTER 1*CLK_P;
DX <= "00000001", "00000010" AFTER 100*CLK_P, "00000001" AFTER 110*CLK_P;
NB <= "00000010", "00000001" AFTER 100*CLK_P, "00000001" AFTER 110*CLK_P;                                   
END control_arch;
